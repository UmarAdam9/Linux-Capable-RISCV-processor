
//=======================================================
//  module declaration
//=======================================================

module m_RISCV32I_ZICSR    import risc_v_core_pkg::* ,tracer_pkg::*;
(
  input                clk_in                ,
  input                rst_in                ,
  
  //MMU interface
  output logic 		  i_req						,		
  output	logic			  i_kill						,			//needed??
  output logic[31:0]	  i_vaddr					,
  output logic			  icache_flush				,
  input 	logic			  i_page_fault				,
  input  logic[31:0]   i_paddr					,
  // i_hit not needed??
  //MMU talks to the instruction cache itself
  
  
  //data bus interface
  input logic[31:0]    dbus_rdata_in			,
  input logic			  dbus_ack_in				,
  
  
  output logic[31:0]  dbus_addr_o				,				//length
  output logic 		 dbus_ld_req_o				,
  output logic 		 dbus_st_req_o				,
  output logic[31:0]  dbus_W_data_o				,				//length
  output logic[3:0]	 dbus_byte_en				,
  
  //also send byte_en??


  
  //mmu interface
  input logic 			  ld_page_fault_in		,
  input logic 			  st_page_fault_in		,
  input logic[31:0] 	  d_paddr_in				,
  input logic 			  d_hit_in					,
  
  	output logic  		 satp_ppn_o					,
	output logic  		 en_vaddr_o					,
	output logic  		 mxr_o						,
	output logic  		 tlb_flush_o				,
	output logic  		 lsu_flush_o				,
	output logic  		 en_ld_st_vaddr_o			,
	output logic  		 dcache_flush_o			,
	output logic  		 sum_o						,
	output logic[1:0]  priv_mode_o				, 				//length??
	output logic[31:0] d_vaddr_o					,
	output logic       d_req_o						,
	output logic       st_req_o
  

	
);

//=======================================================
//  REG/WIRE declarations
//=======================================================

  //Fetch stage 
    //pc + 4 block 
      wire [31:0] PCout_plus4;		
	//pc_mux block				-Umar Adam : commented out the previous mux block
		//wire [31:0] mux_outpc;
	 //pc address						-Umar Adam
		wire [31:0] pc_selector_out;	
	 //exception request wire		-Umar Adam
		wire 			exc_req_if2id;	
	//exception code wire 			-Umar Adam
		wire [3:0]	exc_code_if2id;
    //PC Register block
      wire [31:0] PC_out; 
    //Instruction Memory
      wire [31:0] inst_mem_out;
    //Register
      reg  [31:0] PC_out_reg;
    //Instruction Decoder block
      instruction_t   instruction_o;
		
	 //exception request				-Adam
		wire 			exc_req_out;
	 //exception code					-Adam
		wire [3:0]	exc_code_out;
		

  //Decode stage 
    //hazard detection unit   
		wire			exe_pc_req_fb2if;		//	-Adam
		wire			csr_pc_reqid_fb2if;	//	-Adam
		wire			wfi_req_fb2if;			// -Adam
		wire        PCWrite; 
      wire        IF_DWrite; 
      wire        hazard_out;
    //Register									// why??
      reg         hazard_out_reg; 
      reg         IF_Dwrite_reg;
      reg         PCSrc_reg;
    //PC Register block
      wire [31:0] PC_out_IF_ID; 
    //Instruction Register block
      wire [31:0] inst_out_IF_ID;
    //Register File unit
      wire [31:0] rs1_out; 
      wire [31:0] rs2_out; 
      wire [31:0] rd_regfile;
    //Immediate Generator Block
      wire [31:0] inst_out_imm; 
    //Control Unit 
      wire        RegWrite; 
      wire        MemtoReg; 
      wire        MemRead; 
      wire        MemWrite; 
      wire        jal; 
      wire        jalr;
      wire [1:0]  ALUOp; 
      wire [1:0]  ALUSrcA; 
      wire [1:0]  ALUSrcB;
      wire [5:0]  Branch;
      wire        valid;
		wire [1:0]	csr_ops;					//-Adam
		wire [2:0] 	sys_ops;					//-Adam
		wire			exc_req_out_cntrl;	//-Adam
		wire [3:0]	exc_code_out_cntrl;	//-Adam
    //control_signals_mux block
      wire [33:0] cntrl_out; 				//Umar Adam: change the amount of signals!!!!! [edit: DONE]

		//exception code register block		-Adam
		wire [3:0]	exc_code_out_IF_ID;
	 //exception request	register block		-Adam
		wire 			exc_req_out_IF_ID;
		
		
			
	
		
  //Execute stage 
  
  
	
	
    //PC Register block
      wire [31:0] PC_out_ID_EX; 
    //Instruction Register block
      wire [31:0] inst_out_ID_EX;
    //Immediate Register block 
      wire [31:0] imm_out_ID_EX;
    //Control Signals Register block 	-Umar Adam: change the length to 34 to accomodate the zicsr signals	
      wire [33:0] cntrl_out_ID_EX;
    //rs1 Register block
      wire [31:0] rs1_out_ID_EX;
    //rs2 Register block 
      wire [31:0] rs2_out_ID_EX;
    //jump mux block
      wire [31:0] mux_out_jump;
    //Adder block
      wire [31:0] jump_addr;
    //forwarding unit
      wire [1 :0] forwardA; 
      wire [1 :0] forwardB;
    //rs1 mux block
      wire [31:0] rs1_forwarded;
    //rs2 mux block 
      wire [31:0] rs2_forwarded;
    //ALU_input_A mux block
      wire [31:0] alu_input_A;
    //ALU_input_B mux block
      wire [31:0] alu_input_B;
    //ALU control block
      wire [4 :0] alu_contrl;
    //ALU Block
      wire [31:0] alu_result;
      wire zero; 
      wire nzero; 
      wire less; 
      wire greater; 
      wire lessun; 
      wire greaterun;
    //branch signals
      wire a_n_d_1, a_n_d_2, a_n_d_3, a_n_d_4, a_n_d_5, a_n_d_6;
    //jump signal
      wire PCSrc; 
	 //csr_rw_check block	-Adam
		wire	csr_rd_req;
		wire	csr_wr_req;
		wire	reg_write_exe;
  
  //Memory stage 
    //store unit
      wire [3:0] byte_en;
    //Data memory
      wire [31:0] data_mem_out;
    //control signals Register block
      wire [33:0] cntrl_out_Ex_MEM;
    //ALU Result Register block
      wire [31:0] alu_result_EX_MEM;
    //Instruction Register block
      wire [31:0] inst_out_EX_MEM;
	 //PC register block			-Adam
		logic [31:0] PC_out_EX_MEM;
    //data mem write data mux
      wire [31:0] dmem_wr_data;
    //dmem address selection 
		logic       dmem_addr_sel;
	 //csr_rd_req and csr_wr_req Register blocks
		wire			csr_rd_req_EX_MEM;
		wire			csr_wr_req_EX_MEM;
	 
	 
	 //Csr unit									-Adam
		//fetch[complete signals]
			wire [31:0]	pc_new_csr2if_fb;
			//icache_flush_csr2if_fb??
			//irq_req (for imprecise interrupt handling[will not support])
		//decode[complete signals]
			wire [1:0]  priv_mode_csr2id_fb;
		//WriteBack [complete signals]
			wire [31:0] rdata_csr2wb;	
		//Hazard[complete signals]
			wire 			wfi_req_csr2hzd;
			wire			csr_pc_req_csr2hzd;
			wire			csr_read_req_csr2hzd;
			wire			irq_flush_mem2wb_csr2hzd;
		//LSU	[complete signals]
		   wire [21:0]	satp_ppn_csr2lsu;  //ppn width 22
			wire        en_vaddr_csr2lsu;
			wire			en_ld_st_vaddr_csr2lsu;
			wire			mxr_csr2lsu; 
			wire			lsu_flush_csr2lsu;  
			wire			tlb_flush_csr2lsu;
			wire	      dcache_flush_csr2lsu;
			wire 			sum_csr2lsu;
			wire [1:0]  priv_mode_csr2lsu;  //check length
		
		
		
		//lsu wires		-Adam
			wire dbus_addr_lsu2csr;
			wire ld_page_fault_lsu2csr;
			wire st_page_fault_lsu2csr;
			wire dcache_flush_or_ack_lsu2csr;
		
    
  //Writeback stage 
    //control signals Register block
      wire [23:0] cntrl_out_MEM_WB;
    //data memory Register block
      wire [31:0] dataout_MEM_WB;
    //ALU Result Register block
      wire [31:0] alu_result_MEM_WB;
    //Instruction Register block
      wire [31:0] inst_out_MEM_WB; 
    //Load Unit
      wire [31:0] load_store_unit_out;
    //Writeback mux block
      wire  [31:0]  regfile_write_data; 
      logic [31:0]  regfile_wr_data_final;
    //Instruction Decoder block
      instruction_t   instruction_WB;
  
  //Compression Extension
    wire [31:0] inst_out_comp;
    wire        pc_disable;
	 fsm_state   comp_state;
    wire [31:0] mux_jump_out;
    wire [31:0] dummypc;
    reg  [31:0] dummy_pc_ifid; 
    reg  [31:0] dummy_pc_idex; 
    reg  [31:0] dummy_pc_exmem; 
    reg  [31:0] dummy_pc_memwb;
    reg         compressed; 
    reg         compressed1; 
    reg         compressed2; 
	  
  //atomic extension 
    wire        regfile_rd_addr_sel;
    //wire [1:0]  is_sc_reg_wr;
    wire        dmem_wr_data_sel;
    logic       reserved;
    //amo_controls_t atomic_control_out;
    wire [31:0]   rs2_out_MEM_WB; 
    logic         amo_stall ;
    logic [1:0]   amo_ALUSrcA   ;
    logic [1:0]   amo_ALUSrcB   ;
    logic [1:0]   amo_ALUOp     ;
    logic         amo_MemRead   ;
    logic         amo_MemWrite  ;
    logic         amo_regfile_rd_addr_sel   ;
    logic         amo_RegWrite  ;
    logic         amo_MemtoReg  ;
    logic         amo_dmem_wr_data_sel      ;
    logic [1:0]   amo_is_sc_reg_wr         ;
    logic         is_atomic;
    logic [23:0]  cntrl_out_normal;
    logic         is_atomic_reg;
    logic         is_atomic_reg2;
    logic         is_atomic_reg3;
    logic         amo_stall_reg;
    logic         atomic_;
    logic         lr_w_inst_reg;
    logic         sc_w_inst_reg;
    logic         sc_w_inst_reg2;
    logic         lr_sc_w_inst_reg;
    logic         reserved_reg;
    logic         reserved_reg2;
    logic [31:0]  rs2_forwarded_reg;
    logic         amo_dmem_addr_sel;
    logic         dmem_addr_sel_reg;
    logic         sc_w_inst_EX_MEM;
    logic         sc_w_inst_MEM_WB;
    logic         atomic_stall;
    logic         PCSrc_reg2;
    logic         atomic_stall_2;
//=======================================================
//  Structural Code
//=======================================================

//========================================================================================================
//                                             Fetch Stage
//========================================================================================================
  //(PC + 4) block     OK
    adder pc_adder(
      .a(PC_out     ),
      .b(32'd4      ),
      .c(PCout_plus4)
    );

//  //mux to select (PC + 4) or jump address OK
//    mux mux_pc(
//      .a(PCout_plus4), 
//      .b(jump_addr  ),             
//      .s(PCSrc      ), 
//      .c(mux_outpc  )
//    );
	 
	 
	 //PC selector module   - Umar Adam
	 
	 m_PC_selector selector(
	 	.csr_new_pc_req(csr_pc_reqid_fb2if),
		.exe_new_pc_req(exe_pc_req_fb2if),
		.wfi_req(wfi_req_fb2if),
		.csr_new_pc(pc_new_csr2if_fb),
		.pc_plus_4(PCout_plus4),
		.pc_ff(PC_out),      
		.exe_new_pc(jump_addr),
		.pc_next(pc_selector_out)


	 
	 );
	 
	 
	 
	 
	 
	 
	 

  //PC Register	OK
    register_en   
    #(
      .Default_val(32'h80000000)
    )  PC (  
        .clk  (clk_in                ), 
        .reset(rst_in                ),
        .en   (PCWrite & ~pc_disable & !atomic_stall ),
        .d    ({pc_selector_out[31:1],1'b0}),
        .q    (PC_out                )
    );

  //assigning values to Instruction Memory (FETCH stage) OK 
//    assign mem_ntv_interface_imem.addr     = PC_out;
//    assign mem_ntv_interface_imem.r_en     = PCWrite & ~pc_disable & !atomic_stall ;  
//    assign inst_mem_out                    = mem_ntv_interface_imem.rdata;


	//Assigning values to the MMU interface	-Adam
	assign i_vaddr = PC_out;
// assign i_req	= 1b'1;
	assign i_kill = csr_pc_reqid_fb2if | exe_pc_req_fb2if;
	
	
	//i_kill and i_page_fault assignments??		EDIT: i_page_fault DONE EDIT: i_page_fault DONE
	
	//	Adam : how to assign i_req???
	
	// Adam : how to add read_enable functionality??? {assign mem_ntv_interface_imem.r_en     = PCWrite & ~pc_disable & !atomic_stall ; } do we even need it?
	


  //for synchronisation of PC with Instruction(PC_out-4)  OK
    always@(posedge clk_in or negedge rst_in)
    begin
      if (!rst_in)
          PC_out_reg <= 32'b0;
      else PC_out_reg <= PC_out;        
    end

  //compression unit that converts 16 bit compressed inst into 32 bit inst  OK
    c_controller		compr(					
      .clk            (clk_in         ),
      .reset          (rst_in         ),
      .instruction_in (i_paddr   ),					//from instruction mem
      .PCWrite        (PCWrite        ),
      //.is_atomic      (is_atomic_reg  ),
      .atomic_        (is_atomic        ),
      .amo_stall      (atomic_stall),
      .instruction_out(inst_out_comp  ),
      .pc_disable     (pc_disable     ),
      .compressed     (compressed     ),
      .PCSrc          (PCSrc          ),
      .PC_jump_addr   (jump_addr      ),
      .comp_state     (comp_state     )
	  );
  
  //Dummy_PC Unit (used for compression extension) OK
    dummy_PC dummy_PC_inst(
      .clk          (clk_in           ),
      .reset        (rst_in           ),
      .enable       (!atomic_stall),      //!amo_stall
      .instruction  (i_paddr     ), 			//from instruction mem
      .PCWrite      (PCWrite          ),
      .PCSrc        (PCSrc            ),
      .PC_jump_addr (jump_addr        ),
      .p_state      (comp_state       ),        
      .dummy_pc     (dummypc          )
				  
	);
  assign atomic_stall = (PCSrc_reg) ? 0 : amo_stall;

	//registering dummy pc to be used in further stages  OK
    always@(posedge clk_in or negedge rst_in)
    begin
      if(!rst_in)begin 
        dummy_pc_ifid  <= 32'd0;
        dummy_pc_idex  <= 32'd0;
        dummy_pc_exmem <= 32'd0;
        dummy_pc_memwb <= 32'd0;
        end
      else begin
        dummy_pc_ifid  <= dummypc;
        dummy_pc_idex  <= dummy_pc_ifid;
        dummy_pc_exmem <= dummy_pc_idex;
        dummy_pc_memwb <= dummy_pc_exmem;
        end
    end

  //converting instruction bits into enum for wave display   OK i guess
    Instruction_reg inst_decoder(
      .instruction    (inst_out_comp), 
      .instruction_o  (instruction_o)
    );

  //register PCSrc (jump indication will be used for flush in later stage)    WHY??
    always@(posedge clk_in or negedge rst_in) 
    begin
      if (!rst_in)
           PCSrc_reg <= 1'b0;
      else PCSrc_reg <= PCSrc;
    end
	 
	 
	 
	 
	 //exception gen module 		-Umar Adam
	 m_exc_gen exc_gen(
	 
	.clk(clk_in),
	.rst(rst_in), 
	.instruction(i_paddr),
	.pc(PC_out),
	.csr_new_pc_req(csr_pc_reqid_fb2if), //from the forward stall unit
	.exe_new_pc_req(exe_pc_req_fb2if), //from the forward stall unit
	.wfi_req(wfi_req_fb2if),        //from the forward stall unit
	.if_stall(IF_Dwrite),		//from the forward stall unit
	.i_page_fault(i_page_fault),   //from the MMU
	.exc_req_o(exc_req_out),
	.exc_code_o(exc_code_out)

	 
	 );
	 
	 
	 

//========================================================================================================
//                                            Decode Stage
//========================================================================================================



	//registering exc_req for decode stage -Adam
	register_en #(1)	IF_ID_exc_req(					//Umar Adam:change the register param to 1 bit
		.clk   (clk_in            ), 
      .reset (rst_in            ),
      .flush (PCSrc | PCSrc_reg ), //Umar Adam: how are they using these flushes?? [change these!!]
      .en    (IF_Dwrite_reg     ), 
      .d     (exc_req_out        ),
      .q     (exc_req_out_IF_ID  )
	);
	
	//registering exc_code for decode stage	-Adam
		register_en #(4)	IF_ID_exc_code(					//Umar Adam:change the register param to 4 bits
		.clk   (clk_in            ), 
      .reset (rst_in            ),
      .flush (PCSrc | PCSrc_reg ), //Umar Adam:  [change these!!]
      .en    (IF_Dwrite_reg     ), 
      .d     (exc_code_out        ),
      .q     (exc_code_out_IF_ID  )
	);
	
	
//  //hazard detection (stall of one cycle if hazard detected)
//    hazard_detection_unit hazard_unit(
//      .ID_EX_rd     (inst_out_IF_ID[11:7]), 
//      .IF_ID_rs1    (inst_out_comp[19:15]),  
//      .IF_ID_rs2    (inst_out_comp[24:20]),  
//      .ID_EX_memread(MemRead | (amo_MemRead && lr_w_inst_reg)), 
//      .opcode       (inst_out_comp[6:0]  ),
//      .PCWrite      (PCWrite             ), // signal used to disable PC     
//      .IF_Dwrite    (IF_Dwrite           ), // signal used to disable IF_ID Registers  
//      .hazard_out   (hazard_out          )  // signal used to select 0 as control signals
//  );
//  
  
  
  //Updated hazard detection (stall of one cycle if hazard detected)  -Umar Adam
  m_hazard_detection_unit hazard_unit2(	
	.ID_EX_rd	(inst_out_IF_ID[11:7]), 
	.IF_ID_rs1	(inst_out_comp[19:15]), 
	.IF_ID_rs2	(inst_out_comp[24:20]),
	.ID_EX_memread(MemRead | (amo_MemRead && lr_w_inst_reg)),
	.opcode (inst_out_comp[6:0]  ),
	.exe_pc_req_i(PCSrc),	//PCsrc signal
	.csr_pc_req_i(csr_pc_req_csr2hzd),
	.wfi_req_i(irq_flush_mem2wb_csr2hzd),
	//  input       irq_flush_mem2wb,
	.exe_pc_req_o(exe_pc_req_fb2if),
	.csr_pc_req_o(csr_pc_reqid_fb2if),
	.wfi_req_o(wfi_req_fb2if),
	.PCWrite(PCWrite), 	 //Blocks the pc read 
	.IF_Dwrite(IF_Dwrite),   //blocks the IF/ID pipeline
	.hazard_out(hazard_out)	 //sends all zeroes as control signals to the execute stage (NOOP?)
  );
  
  
  
  //registering Hazard out and IF_D write 
    always@(posedge clk_in or negedge rst_in)
    begin
      if (!rst_in) begin
          hazard_out_reg <= 1'b0;
          IF_Dwrite_reg  <= 1'b0;
          PCSrc_reg2     <= 0;
      end
      else begin
        hazard_out_reg <= hazard_out;
        IF_Dwrite_reg  <= IF_Dwrite;
        PCSrc_reg2     <= PCSrc_reg;
      end
    end

  //Registering PC For Decode Stage
    register_en IF_ID_pcout(
      .clk   (clk_in            ), 
      .reset (rst_in            ),
      .flush (PCSrc | PCSrc_reg ), //generate flush for two cycle  [Umar Adam: Figure out why 2 flushes!]
      .en    (IF_Dwrite_reg     ), 
      .d     (PC_out_reg        ),
      .q     (PC_out_IF_ID      )
    );

  //Registering Instruction For Decode Stage
    register_en IF_ID_instout(
      .clk   (clk_in            ), 
      .reset (rst_in            ), 
      .flush (PCSrc | PCSrc_reg ), //generate flush for two cycle	[Umar Adam: Figure out why 2 flushes!]
      .en    (IF_Dwrite_reg  & atomic_stall_2  ),  
      .d     (inst_out_comp     ),
      .q     (inst_out_IF_ID    )
    );
    assign atomic_stall_2 = (PCSrc_reg2) ? 1:!amo_stall_reg;
  //mux at input of rd of regfile to select between rd and rs2_out for amo swap instruction
    mux mux_rd_regfile(
      .a(inst_out_MEM_WB[11:7]),    //rd
      .b(inst_out_MEM_WB[24:20]),   //rs2
      .s(cntrl_out_MEM_WB[22]),    //regfile_rd_addr_sel
      .c(rd_regfile)
    );
  //Register File
    register_file reg_file(
      .write_data (regfile_wr_data_final ), 
      .rs1        (inst_out_IF_ID[19:15] ),  
      .rs2        (inst_out_IF_ID[24:20] ),   
      .rd         (inst_out_MEM_WB[11:7] ),     
      .we         (cntrl_out_MEM_WB[1]   ),   //regwrite
      .clk        (clk_in                ), 
      .rst        (rst_in                ),
      .read_data1 (rs1_out               ), 
      .read_data2 (rs2_out               )
  );

  //Immediate Generator
    Imm_Gen imm_gen(
      .Inst_In    (inst_out_IF_ID        ),      
      .Imm_Out    (inst_out_imm          )
  );

//  //Generate control Signals
//    control_unit control_unit(
//      .Op         (inst_out_IF_ID[6:0]   ),              
//      .funct3     (inst_out_IF_ID[14:12] ),        
//      .funct7     (inst_out_IF_ID[31:25] ),
//      .ALUOp      (ALUOp                 ), 
//      .ALUSrcA    (ALUSrcA               ), 
//      .ALUSrcB    (ALUSrcB               ),
//      .Branch     (Branch                ),
//      .RegWrite   (RegWrite              ), 
//      .MemtoReg   (MemtoReg              ), 
//      .MemRead    (MemRead               ), 
//      .MemWrite   (MemWrite              ),
//      .jal        (jal                   ), 
//      .jalr       (jalr                  ),
//      .valid      (valid                 ),
//      .dmem_addr_sel(dmem_addr_sel)
//  );
//  
  
  
  //updated control signals					-Umar Adam
  m_control_unit_ZICSR control_unit2(
  .Op(inst_out_IF_ID[6:0]   ),
  .funct3(inst_out_IF_ID[14:12] ),
  .funct7(inst_out_IF_ID[31:25] ),
  .funct5(inst_out_IF_ID[31:25] ),		//Umar Adam: CHANGE THIS!!!!
  .priv_mode(),
  .ALUOp (ALUOp                 ), 
  .ALUSrcA (ALUSrcA               ), 
  .ALUSrcB(ALUSrcB               ),
  .Branch(Branch                ),
  .RegWrite(RegWrite              ), 
  .MemtoReg(MemtoReg              ), 
  .MemRead(MemRead               ), 
  .MemWrite(MemWrite              ), 
  .jal (jal                   ),
  .jalr(jalr                  ), 
  .valid(valid                 ),
  .dmem_addr_sel(dmem_addr_sel),               //select between alu_out and alu_out_reg
  
  .exc_req_if2id(exc_req_out_IF_ID),				/**Umar Adam : extra signals for zicsr extension**/
  .exc_code_if_id(exc_code_out_IF_ID),
  
  .csr_ops(csr_ops),
  .sys_ops(sys_ops),
  
  .exc_req(exc_req_out_cntrl),
  .exc_code(exc_code_out_cntrl)
 
);
    
  //atomic instructions control unit
    amo_control_unit amo_control_unit_inst(
        .clk(clk_in),
        .reset(rst_in),
        .instruction(inst_out_comp),  //instruction will come from fetch stage 
        //.Instruction_reg(inst_out_IF_ID),
        .lr_sc_w_inst(lr_sc_w_inst),
        .is_atomic(is_atomic),
        .atomic_(atomic_),
        .lr_w_inst_reg(lr_w_inst_reg),
        .sc_w_inst_reg(sc_w_inst_reg),
        .amo_stall(amo_stall),
        .ALUSrcA(amo_ALUSrcA),
        .ALUSrcB(amo_ALUSrcB),  
        .ALUOp(amo_ALUOp),   
        .MemRead(amo_MemRead),
        .MemWrite(amo_MemWrite),
        .regfile_rd_addr_sel(amo_regfile_rd_addr_sel),  
        .RegWrite(amo_RegWrite),
        .MemtoReg(amo_MemtoReg),
        .dmem_wr_data_sel(amo_dmem_wr_data_sel),  
        .dmem_addr_sel(amo_dmem_addr_sel),  
        .is_sc_reg_wr(amo_is_sc_reg_wr)

    );


  //mux to select control signals (18'b0 if there is a stall or flush)
    mux #(34) control_signals(						//Umar Adam : change the mux param to 34 bits and add the zicsr signals [edit:DONE]
      .a({csr_ops[1:0],sys_ops[2:0],exc_req_out_cntrl,exc_code_out_cntrl[3:0],dmem_addr_sel,amo_regfile_rd_addr_sel,amo_stall,amo_is_sc_reg_wr[1:0],amo_dmem_wr_data_sel,ALUOp[1:0], ALUSrcA[1:0], ALUSrcB[1:0], jalr, Branch[5:0], jal, MemRead, MemWrite, RegWrite, MemtoReg }), 
      .b(34'd0), 
      .s(hazard_out_reg | PCSrc), 
      .c(cntrl_out_normal)
  );

  //registering stall signals 
    always_ff @(posedge clk_in or negedge rst_in) begin
      if(!rst_in) begin
        is_atomic_reg <= 0;
        lr_sc_w_inst_reg  <= 0;
        amo_stall_reg <= 0;
        dmem_addr_sel_reg <= 0;
        is_atomic_reg2    <= 0;
        is_atomic_reg3    <= 0;
      end
      else begin 
        is_atomic_reg <= is_atomic;
        amo_stall_reg <= amo_stall;
        lr_sc_w_inst_reg <= lr_sc_w_inst;
        dmem_addr_sel_reg <=  dmem_addr_sel;
        is_atomic_reg2  <= is_atomic_reg;
        is_atomic_reg3    <= is_atomic_reg2;
      end 
    end
  //selecting control signals between atomic controls and normal controls [Umar Adam : Should the zicsr control signals be changed because of atomic controls???]
    mux #(34) final_controls(
      .a(cntrl_out_normal),
      .b({csr_ops[1:0],sys_ops[2:0],exc_req_out_cntrl,exc_code_out_cntrl[3:0],amo_dmem_addr_sel,amo_regfile_rd_addr_sel,amo_stall,amo_is_sc_reg_wr[1:0],amo_dmem_wr_data_sel,amo_ALUOp[1:0], amo_ALUSrcA[1:0],amo_ALUSrcB[1:0],jalr,Branch[5:0],jal,amo_MemRead,amo_MemWrite,amo_RegWrite,amo_MemtoReg}),
      .s(is_atomic_reg | cntrl_out_ID_EX[21] | lr_sc_w_inst_reg),
      .c(cntrl_out)
    );

    //amo_memtoreg = cntrl_out[0]
    //amo_regwrite = cntrl_out[1]
    //amo_memwrite = cntrl_out[2]
    //amo_memread = cntrl_out[3]
    //jal = cntrl_out[4]
    //branch[5:0] = cntrl_out[10:5]
    //jalr = cntrl_out[11]
    //alusrc_b[1:0] = cntrl_out[13:12]
    //alusrc_a[1:0] = cntrl_out[15:14]
    //alu_op[1:0] = cntrl_out[17:16]
    //dmem_wr_dta_sel = cntrl_out[18]
    //is_sc_reg_wr_sel = cntrl_out[20:19]
    //amo_stall = cntrl_out[21]
    //amo_regfile_rd_addr_sel = cntrl_out[22]
    //amo_dmem_addr_sel       = cntrl_out[23]

//========================================================================================================
//                                          Execute Stage
//========================================================================================================



  //Registering PC For Execute Stage
    register ID_EX_pcout(
      .clk   (clk_in                ), 
      .reset (rst_in                ),
      .flush (PCSrc |hazard_out_reg ),   //Umar Adam: why is hazard_out_reg being used??
      .d     (PC_out_IF_ID          ), 
      .q     (PC_out_ID_EX          )
    );

  //Registering Instruction For Execute Stage
    register ID_EX_instout(
      .clk   (clk_in                ), 
      .reset (rst_in                ), 
      .flush (PCSrc |hazard_out_reg ),        //Umar Adam: why is hazard_out_reg being used?? 
      .d     (inst_out_IF_ID        ),   
      .q     (inst_out_ID_EX        )
    );

  //Registering Immediate For Execute Stage
    register ID_EX_imm(
      .clk   (clk_in                ), 
      .reset (rst_in                ), 
      .flush (PCSrc                 ), 
      .d     (inst_out_imm          ), 
      .q     (imm_out_ID_EX         )
    );

  //Registering Controls Signals For Execute Stage		[Umar Adam: changed the length to 34]
    register #(34) ID_EX_controls(
      .clk   (clk_in                ), 
      .reset (rst_in                ), 
      .flush (PCSrc                 ), 
      .d     (cntrl_out             ),
      .q     (cntrl_out_ID_EX       )
    );

  //Registering Rs1_out For Execute Stage
    register ID_EX_rs1out(
      .clk   (clk_in                ), 
      .reset (rst_in                ), 
      .flush (PCSrc                 ), 
      .d     (rs1_out               ), 
      .q     (rs1_out_ID_EX         )
    );

  //Registering Rs2_out For Execute Stage
    register ID_EX_rs2out(
      .clk   (clk_in                ), 
      .reset (rst_in                ), 
      .flush (PCSrc                 ), 
      .d     (rs2_out               ), 
      .q     (rs2_out_ID_EX         )
    );
	 
	 
	 
	 
	 
	 

  //mux that selects rs1 for Jalr or PC for other jumps
    mux jump(
      .a     (dummy_pc_idex         ), 
      .b     (rs1_forwarded         ),   
      .s     (cntrl_out_ID_EX[11]   ), //JALR  
      .c     (mux_out_jump          )
    );

  //adder to calculate jump address for PC
    adder ADDJump_imm(
      .a     (mux_out_jump          ),
      .b     (imm_out_ID_EX         ),
      .c     (jump_addr             )
    );

  //Generate Select lines for mux A and mux B from where to forward data(of rs1 and rs2)
    forwarding_unit forwarding_unit(
      .rs1            (inst_out_ID_EX[19:15]), 
      .rs2            (inst_out_ID_EX[24:20]), 
      .EX_MEM_rd      (inst_out_EX_MEM[11:7]), 
      .MEM_WB_rd      (inst_out_MEM_WB[11:7]),
      .EX_MEM_regwrite(cntrl_out_Ex_MEM[1]  ),  //regwrite
      .MEM_WB_regwrite(cntrl_out_MEM_WB[1]  ),  //regwrite
      .is_atomic      (is_atomic_reg3       ),
      .sc_w_inst_EX_MEM(sc_w_inst_EX_MEM    ),
      .sc_w_inst_MEM_WB(sc_w_inst_MEM_WB    ),
      .reserved       (reserved             ),
      .forward_A      (forwardA             ), 
      .forward_B      (forwardB             )
    );

  //mux to select latest rs1 data using forwarding 
    mux_4x1 mux_rs1(
      .a     (rs1_out_ID_EX         ),  
      .b     (regfile_write_data    ), //mem hazard   
      .c     (alu_result_EX_MEM     ), //execute hazard
      .d     ((reserved_reg) ? 0:1  ),  //when sc.w hazard occurs this will go 
      .s     (forwardA              ), 
      .q     (rs1_forwarded         )
    );

  //mux to select latest rs2 data using forwarding 
    mux_4x1 mux_rs2(
      .a     (rs2_out_ID_EX         ),  
      .b     (regfile_write_data    ), //mem hazard  
      .c     (alu_result_EX_MEM     ), //execute hazard
      .d     ((reserved_reg) ? 0:1  ),
      .s     (forwardB              ),  
      .q     (rs2_forwarded         )
    );

  //registering compressed signal from fetch stage to be used in execute
	  always@(posedge clk_in or negedge rst_in)			
	  begin
      if(!rst_in)begin 
          compressed1       <= 1'b0;
          compressed2       <= 1'b0;
          sc_w_inst_reg2    <= 0;  
          sc_w_inst_EX_MEM  <= 0;    
          sc_w_inst_MEM_WB  <= 0;
      end
      else begin
          compressed1       <= compressed;
          compressed2       <= compressed1;
          sc_w_inst_reg2    <= sc_w_inst_reg;      //this is in execute stage now
          sc_w_inst_EX_MEM  <= sc_w_inst_reg2;   //this is in memory stage now
          sc_w_inst_MEM_WB  <= sc_w_inst_EX_MEM; //this is in write back stage now
      end
	  end

  //mux to select "2" (rd=pc+2) when there is compressed instruction
	  mux comp_jump (
      .a	(32'd4          ),
      .b	(32'd2          ), 
      .s	(compressed2    ), 
      .c	(mux_jump_out   )
	  );

  //mux to select input For ALU First(A) input
    mux_4x1 mux_ALU_A(
      .a     (rs1_forwarded         ), 
      .b     (dummy_pc_idex         ), 
      .c     (32'd0                 ),
      .d     (data_mem_out          ),  //comes directly from main memory 
      .s     (cntrl_out_ID_EX[15:14]),  //ALUSrcA
      .q     (alu_input_A           )
    );
  
  //mux to select input For ALU Second(B) input
    mux_4x1 mux_ALU_B(
      .a     (rs2_forwarded         ), 
      .b     (imm_out_ID_EX         ), 
      .c     (mux_jump_out          ),
      .d     (32'd0                 ),    //for atomic rs1+0 to get M[rs1]         
      .s     (cntrl_out_ID_EX[13:12]),  //ALUSrcB
      .q     (alu_input_B           )
    );

  //Generate control lines for ALU 
    ALUControl alu_control(
      .ALUOp          (cntrl_out_ID_EX[17:16]), 
      .funct3         (inst_out_ID_EX[14:12] ), 
      .funct7         (inst_out_ID_EX[31:25] ),
      .funct5         (inst_out_ID_EX[31:27] ),   
      .OP             (inst_out_ID_EX[6:0]   ),
      .ALUCtl         (alu_contrl            )
    );

  //ALU Unit
    ALU alu (
      .ALUctl         (alu_contrl            ), 
      .A              (alu_input_A           ), 
      .B              (alu_input_B           ), 
      .ALUOut         (alu_result            ), 
      .Zero           (zero                  ),
      .n_zero         (nzero                 ),
      .less_than      (less                  ),
      .greater_than   (greater               ),
      .less_than_u    (lessun                ),
      .greater_than_u (greaterun             )
    );
	 
	 
	 //csr_rw_checker module 	-Umar Adam
	 
	 m_csr_RWChecker csr_rw_checker(

		.instruction(inst_out_ID_EX), 	
		.immediate(imm_out_ID_EX), 		
		.csr_ops(cntrl_out_ID_EX[33:32]),
		.RegWrite_id2exe(cntrl_out_ID_EX[1]),

		.csr_rd_req(csr_rd_req),
		.csr_wr_req(csr_wr_req),
		.RegWrite(reg_write_exe) 		//Register this RegWrite signal for the next pipeline stage 

);
	 
	 
	 

  //Checking different Branch Conditions
    assign a_n_d_1 = zero       & cntrl_out_ID_EX[5]; //BEQ
    assign a_n_d_2 = nzero      & cntrl_out_ID_EX[6]; //BNE
    assign a_n_d_3 = less       & cntrl_out_ID_EX[7]; //BLT
    assign a_n_d_4 = greater    & cntrl_out_ID_EX[8]; //BGE
    assign a_n_d_5 = lessun     & cntrl_out_ID_EX[9]; //BLTU
    assign a_n_d_6 = greaterun  & cntrl_out_ID_EX[10];//BGEU

  //PCSRC is 1 if any of Jump condition is true (Branch , Jalr or Jal)
    assign PCSrc = a_n_d_1 | a_n_d_2 |a_n_d_3 |a_n_d_4 |a_n_d_5 |a_n_d_6 | cntrl_out_ID_EX[11] | cntrl_out_ID_EX[4];


//========================================================================================================
//                                         Memory Stage
//========================================================================================================

  // Generate byte_enable for data memory		//UA : Okay
    store_unit store_unit(
      .func3       (inst_out_ID_EX[14:12] ),
      .dmem_address(alu_result[1:0]       ), 
      .byte_en     (byte_en               )
    );

  //registering rs2 forwarded										EDIT: UA: WHYY???
  always_ff @(posedge clk_in or negedge rst_in) begin
    if(!rst_in)
      rs2_forwarded_reg <= 0;
    else  
      rs2_forwarded_reg <= rs2_forwarded;
  end
 


 //mux that selects the data to be written in data memory {Umar Adam: NEW EDIT: for AMO instructions}
    mux dmem_wr_mux(
      .a(rs2_forwarded), //rs2_forwarded_reg
      .b(alu_result),
      .s(cntrl_out_ID_EX[18]),  //amo_dmem_wr_data_sel
      .c(dmem_wr_data)
    );
	 
	 
	 
	 
	 
  // Assigning values to Data Memory
  // Sending unregistered values(execute stage) to Data Memory because our memory is input registered
   /*  assign mem_ntv_interface_dmem.addr        = (cntrl_out_ID_EX[23]) ? alu_result : alu_result_EX_MEM;   //amo_dmem_addr_sel      
    assign mem_ntv_interface_dmem.wdata       = dmem_wr_data;             
    assign mem_ntv_interface_dmem.w_en        = reserved | cntrl_out_ID_EX[2];   
    assign mem_ntv_interface_dmem.r_en        = cntrl_out_ID_EX[3];   
    assign mem_ntv_interface_dmem.byteenable  = byte_en;
    assign data_mem_out                       = mem_ntv_interface_dmem.rdata; */



  //atomic reservation file for lr.w/sc.w instructions 
    reservation_file  reserve_file(
          .clk(clk_in),
          .rst(rst_in),
          .instruction(inst_out_ID_EX),
          .reserved(reserved)
    );


  //Registering Controls Signals For Memory Stage  [Umar Adam:why is the register 23 and not 24? also changed it to 34]
    register #(34) EX_MEM_controls(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     ({cntrl_out_ID_EX[33:2],reg_write_exe ,cntrl_out_ID_EX[0]} ),
      .q     (cntrl_out_Ex_MEM     )
    );
	 

  //Registering ALU Result For Memory Stage
    register EX_MEM_ALU(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     (alu_result           ), 
      .q     (alu_result_EX_MEM    )
    );

  //Registering Instruction For Memory Stage
    register EX_MEM_instout(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     (inst_out_ID_EX       ), 
      .q     (inst_out_EX_MEM      )
    );
	 
	 
	 //register csr_rd_req and wr_req for csr module    -Umar Adam 
	 register #(1) EX_MEM_csr_rd_req(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     (csr_rd_req      ), 
      .q     (csr_rd_req_EX_MEM      )
    );
	 

	 register #(1) EX_MEM_csr_wr_req(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     (csr_wr_req      ), 
      .q     (csr_wr_req_EX_MEM      )
		
    );
	 
	 
	 
	 
	 
	 //register fence_i req (first generate it lol)
	 
	 
	 
	 //register PC						
	  register EX_MEM_pcout(
      .clk   (clk_in                ), 
      .reset (rst_in                ),											
      .d     (PC_out_ID_EX          ), 
      .q     (PC_out_EX_MEM)
    );
	 
	 
	 
	 
	 //instantiate the LSU module		-Adam
	 
	 m_lsu lsu(			
	
		.alu_result((cntrl_out_ID_EX[23]) ? alu_result : alu_result_EX_MEM),
		.write_data(dmem_wr_data),
		.mem_rd(cntrl_out_ID_EX[3]),
		.mem_wr(reserved | cntrl_out_ID_EX[2]),
		.byte_enable_in(byte_en),
		
		.satp_ppn(satp_ppn_csr2lsu),
		.en_vaddr(en_vaddr_csr2lsu),
		.mxr(mxr_csr2lsu),
		.tlb_flush(tlb_flush_csr2lsu),
		.en_ld_st_vaddr(en_ld_st_vaddr_csr2lsu),
		.dcache_flush(dcache_flush_csr2lsu),
		.sum(sum_csr2lsu),
		.priv_mode(priv_mode_csr2lsu),
		
		.dbus_rdata(dbus_rdata_in),
		.dbus_ack(dbus_ack_in),
		
		
		.ld_page_fault(ld_page_fault_in),
		.st_page_fault(st_page_fault_in),
		.d_paddr(d_paddr_in),
		.d_hit(d_hit_in),
		
		.hzd2lsu_lsu_flush('0),   //from hazard unit
		
		.lsu2csr_dbus_addr(dbus_addr_lsu2csr),
		.lsu2csr_ld_page_fault(ld_page_fault_lsu2csr),
		.lsu2csr_st_page_fault(st_page_fault_lsu2csr),
		.lsu2csr_dcache_flush_or_ack(dcache_flush_or_ack_lsu2csr),
		
		.lsu_req(),					//To hazard unit  (These stalls are yet to be implemented btw)
		.lsu_ack(),
		
		.r_data(),				//To WB stage
		
		.lsu2mmu_satp_ppn(satp_ppn_o),	//To mmu outside the core
		.lsu2mmu_en_vaddr(en_vaddr_o),
		.lsu2mmu_mxr(mxr_o),
		.lsu2mmu_tlb_flush(tlb_flush_o),
		.lsu2mmu_lsu_flush(lsu_flush_o),
		.lsu2mmu_en_ld_st_vaddr(en_ld_st_vaddr_o),
		.lsu2mmu_dcache_flush(dcache_flush_o),
		.lsu2mmu_sum(sum_o),
		.lsu2mmu_priv_mode(priv_mode_o),
		.lsu2mmu_d_vaddr(d_vaddr_o),
		.lsu2mmu_d_req(d_req_o),
		.lsu2mmu_st_req(st_req_o),
		
									
		.dbus_addr(dbus_addr_o),						//To data bus outside the core
		.lsu2dbus_ld_req(dbus_ld_req_o),
		.lsu2dbus_byte_enable(dbus_byte_en),
		.lsu2dbus_st_req(dbus_st_req_o),
		.lsu2dbus_W_data(dbus_W_data_o)

	 
	 );
	 
	 
	 
	 
	 //instantiating the csr module
	 
	 m_csr_new csr(
	 
		.rst(rst_in),
		.clk(clk_in),


		//inputs from other units ===========================

		//EXECUTE unit <---> CSR  
		.csr_ops_in(cntrl_out_Ex_MEM[33:32]),			//check the width
		.sys_ops_in(cntrl_out_Ex_MEM[31:29]),			//check the width
		.exc_req_in(cntrl_out_Ex_MEM[28]),
		.irq_req_in('0),
		.csr_rd_req_in(csr_rd_req_EX_MEM),
		.csr_wr_req_in(csr_wr_req_EX_MEM),
		.fence_i_req_in('0),    					//not implemented yet

		.csr_addr_in(inst_out_EX_MEM[31:20]),		//check the length , comes from the instruction
		.pc_in(PC_out_EX_MEM),
		.instr_in(inst_out_EX_MEM),
		.csr_wdata_in(alu_result_EX_MEM),     //comes from the ALU
		.exc_code_in(cntrl_out_Ex_MEM[27:24]),		//check the length
		.instr_flushed_in(),

		//HZD <---> CSR unit 
		.pipe_stall_in('0),			//comes from lsu_div_stall which is yet to be implemented

		//CLINT <---> CSR 
		.timer_val_low_in('0), 
		.timer_val_high_in('0),  

		//SOC <---> CSR  
		.csr_mhartid_in('0),                           
		.ext_irq_in('0),  
		.timer_irq_in('0),  
		.soft_irq_in('0),
		.uart_irq_in('0),   

		//LSU <---> CSR 
		.dbus_addr_in(dbus_addr_lsu2csr),
		.ld_page_fault_in(ld_page_fault_lsu2csr),
		.st_page_fault_in(st_page_fault_lsu2csr),
		.pc_next_in('0),
		.dcache_flush_ack_in(dcache_flush_or_ack_lsu2csr),
		//outputs to other units===========================

		//CSR <---> WRITE_BACK  
		.csr_rdata_o(rdata_csr2wb),  

		//CSR <---> HZD
		.new_pc_req_o(csr_pc_req_csr2hzd), 
		.irq_flush_lsu_o(irq_flush_mem2wb_csr2hzd),
		.wfi_req_o(wfi_req_csr2hzd ),
		.csr_read_req_o(csr_read_req_csr2hzd),
		
		//CSR <---> DECODE unit feedback 
		.priv_mode_o(priv_mode_csr2id_fb),

		//CSR <---> FETCH unit feedback
		.pc_new_o(pc_new_csr2if_fb),	
		.icache_flush_o(icache_flush),

		//CSR <---> LSU unit
		.satp_ppn(satp_ppn_csr2lsu),  //is the width correct????
		.en_vaddr(en_vaddr_csr2lsu),
		.mxr(mxr_csr2lsu),
		.tlb_flush(tlb_flush_csr2lsu),
		.en_ld_st_vaddr(en_ld_st_vaddr_csr2lsu),
		.dcache_flush(dcache_flush_csr2lsu),
		.sum(sum_csr2lsu),
		.priv_mode_to_lsu(priv_mode_csr2lsu),
		.lsu_flush(),//useless??
		
		
		
		
		//debug
		.mcause_o(),
		.mepc_o(),
		.mtval_o()

		
			 
			 
	 
	 
	 );
	 
	 
	 
	 
	 
	 
	 
	 

//========================================================================================================
//                                         Writeback Stage
//========================================================================================================

  //Registering Controls Signals For Writeback Stage
    register #(23) MEM_WB_controls(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     (cntrl_out_Ex_MEM),
      .q     (cntrl_out_MEM_WB     )
    );

  //Registering Datamemory Out For Writeback Stage
    register MEM_WB_datamem(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     (data_mem_out         ), 	//take care of data_mem_out -Adam
      .q     (dataout_MEM_WB       )
    );
  
  //Registering ALU Result for Writeback Stage
    register MEM_WB_ALU(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     (alu_result_EX_MEM    ), 
      .q     (alu_result_MEM_WB    )
    );

  //Registering Instruction for Writeback Stage
    register MEM_WB_instout(
      .clk   (clk_in               ), 
      .reset (rst_in               ), 
      .d     (inst_out_EX_MEM      ), 
      .q     (inst_out_MEM_WB      )
    );
  
  //Generates data to be loaded in Register file for load instruction
    load_unit load_unit(
      .data_in_load (dataout_MEM_WB        ), 
      .func3        (inst_out_MEM_WB[14:12]),  
      .addr         (alu_result_MEM_WB[1:0]),  
      .data_out_load(load_store_unit_out   )
    );

  //Selects data to be written in register file (load_unit_out or Alu_result)
    mux write_back(
      .a     (alu_result_MEM_WB    ),  
      .b     (load_store_unit_out  ),  
      .s     (cntrl_out_MEM_WB[0]  ), //memtoreg
      .c     (regfile_write_data   )
    );

  //registering reserved signal
    always_ff @(posedge clk_in or negedge rst_in) begin
      if(!rst_in) begin 
        reserved_reg <= 0;
        reserved_reg2 <= 0;
        end
      else begin 
        reserved_reg <= reserved; 
        reserved_reg2 <= reserved_reg;
        end
      end

    //final selection for data to be written in register file 
    mux_4x1 final_write_back(
      .a(regfile_write_data),       //in case of no sc.w instruction
      .b((reserved_reg2) ? 32'd0: 32'd1),                    //in case of sc.w success
      .c(32'd1),                    //in case of sc.w failure
      .d(rs2_out_MEM_WB),
      .s(cntrl_out_MEM_WB[20:19]), // is_sc_reg_write
      .q(regfile_wr_data_final)                          //mux out
    );
	 
	 
  //converting instruction bits into enum for wave display
    Instruction_reg inst_decoder_WB(
      .instruction    (inst_out_MEM_WB ), 
      .instruction_o  (instruction_WB)
    );


endmodule
